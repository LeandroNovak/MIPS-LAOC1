LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY control IS
	PORT(
		Opcode			:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		clock, reset	:IN STD_LOGIC;
		RegDst			:OUT STD_LOGIC;
		ALUSrc			:OUT STD_LOGIC;
		MemtoReg			:OUT STD_LOGIC;
		RegWritej		:OUT STD_LOGIC;
		MemRead			:OUT STD_LOGIC;
		Branch			:OUT STD_LOGIC;
		ALUop				:OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END control;

ARCHITECTURE behavior OF control IS
	SIGNAL R_format, Lw, Sw, Beq :STD_LOGIC;
BEGIN
	R_format		<='1' WHEN Opcode ="000000" ELSE '0';
	Lw				<='1' WHEN Opcode ="100011" ELSE '0';
	Sw				<='1' WHEN Opcode ="101011" ELSE '0';
	Beq			<='1' WHEN Opcode ="000100" ELSE '0';

	RegDst		<=R_format;
	ALUSrc		<=Lw OR Sw;
	MemtoReg		<=Lw;
	RegWritej	<=R_format OR Lw;
	MemRead		<=Lw;
	Branch		<=Beq;
	ALUop(1)		<=R_format;
	ALUop(0)		<=Beq;
END behavior;